`include "environment.sv"

program test(intf vif);
    bit read;
	bit write;
 	environment env;
 	task test1();
    // 	env.gen.INCR4(write);
	endtask

    initial begin
    end

endprogram