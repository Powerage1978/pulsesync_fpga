`timescale 1ns / 1ps

package sys_pkg;
    parameter C_SYS_FREQ = 32'd50000000;   // 50 MHz
endpackage