`timescale 1ns / 1ps

package sim_pkg;
    parameter C_CLOCK_PERIOD = 20;
    parameter C_HALF_PERIOD = C_CLOCK_PERIOD / 2;
endpackage