`timescale 1ns / 1ps

package gatedriver_pkg;
    parameter C_COUNT_SIZE = 25;
    parameter C_IDX_SIZE = 4;
    parameter C_OUTPUT_WIDTH = 4;
    parameter C_WORD_SIZE = 32;
    parameter C_NO_OF_STATES_OFFSET = 8;
    parameter C_T_TOLERANCE = 100;
    parameter C_STATUS_SIZE = 3;
endpackage