`timescale 1ns / 100ps

/*
 * Defines system wide parameters.
 */
package sys_pkg;
    parameter C_SYS_FREQ = 32'd50000000;   // 50 MHz logic frequency, must match settings definied within Vivado project
endpackage